`timescale 1ns / 10ps

module cordic_17(in, iout, qout, ain, clk);
   input [19:0]    ain;
   input [16:0]    in;
   output [16:0]   iout, qout;
   input           clk;
   reg [18:0]     a0;
   reg [17:0]     a1;
   reg [17:0]     a2;
   reg [16:0]     a3;
   reg [15:0]     a4;
   reg [14:0]     a5;
   reg [13:0]     a6;
   reg [12:0]     a7;
   reg [11:0]     a8;
   reg [10:0]     a9;
   reg [9:0]      a10;
   reg [8:0]      a11;
   reg [7:0]      a12;
   reg [6:0]      a13;
   reg [5:0]      a14;
   reg [4:0]      a15;
   reg [16:0]     i1, i2, i3, i4, i5, i6, i7, i8, i9;
   reg [16:0]     i10, i11, i12, i13, i14, i15, i16, i17;
   reg [16:0]     q0, q1, q2, q3, q4, q5, q6, q7, q8, q9;
   reg [16:0]     q10, q11, q12, q13, q14, q15, q16, q17;
   always @ (posedge clk)
     begin
        /* 90 degrees */
        a0[17:0]  <= ain[17:0];
        a0[18] <= ~ain[18];
        if(ain[19])
          q0 <= -in;
        else
          q0 <= in;
        /* 45 degrees */
        a1[16:0] <= a0[16:0];
        a1[17] <= ~a0[17];
        q1 <= q0;
        q1 <= q0;
        if(a0[18])
          i1 <= q0;
        else
          i1 <= -q0;
        /* 26.56 degrees */
        if(a1[17])
          begin
             a2 <= a1 + 18'd77376;
             i2 <= i1 + {q1[16], q1[16:1]};
             q2 <= q1 - {i1[16], i1[16:1]};
          end
        else
          begin
             a2 <= a1 - 18'd77376;
             i2 <= i1 - {q1[16], q1[16:1]};
             q2 <= q1 + {i1[16], i1[16:1]};
          end // else: !if(a1[17])
        /* 14.036 degrees */
        if(a2[17])
          begin
             a3 <= a2[16:0] + 17'd40884;
             i3 <= i2 + {{2{q2[16]}}, q2[16:2]};
             q3 <= q2 - {{2{i2[16]}}, i2[16:2]};
          end
        else
          begin
             a3 <= a2[16:0] - 17'd40884;
             i3 <= i2 - {{2{q2[16]}}, q2[16:2]};
             q3 <= q2 + {{2{i2[16]}}, i2[16:2]};
          end // else: !if(a2[17])
        /* 7.125 degrees */
        if(a3[16])
          begin
             a4 <= a3[15:0] + 16'd20753;
             i4 <= i3 + {{3{q3[16]}}, q3[16:3]};
             q4 <= q3 - {{3{i3[16]}}, i3[16:3]};
          end
        else
          begin
             a4 <= a3[15:0] - 16'd20753;
             i4 <= i3 - {{3{q3[16]}}, q3[16:3]};
             q4 <= q3 + {{3{i3[16]}}, i3[16:3]};
          end // else: !if(a3[16])
        /* 3.576 degrees */
        if(a4[15])
          begin
             a5 <= a4[14:0] + 15'd10417;
             i5 <= i4 + {{4{q4[16]}}, q4[16:4]};
             q5 <= q4 - {{4{i4[16]}}, i4[16:4]};
          end
        else
          begin
             a5 <= a4[14:0] - 15'd10417;
             i5 <= i4 - {{4{q4[16]}}, q4[16:4]};
             q5 <= q4 + {{4{i4[16]}}, i4[16:4]};
          end // else: !if(a4[15])
        /* 1.790 degrees */
        if(a5[14])
          begin
             a6 <= a5[13:0] + 14'd5213;
             i6 <= i5 + {{5{q5[16]}}, q5[16:5]};
             q6 <= q5 - {{5{i5[16]}}, i5[16:5]};
          end
        else
          begin
             a6 <= a5[13:0] - 14'd5213;
             i6 <= i5 - {{5{q5[16]}}, q5[16:5]};
             q6 <= q5 + {{5{i5[16]}}, i5[16:5]};
          end // else: !if(a5[14])
        /* 0.895 degrees */
        if(a6[13])
          begin
             a7 <= a6[12:0] + 13'd2607;
             i7 <= i6 + {{6{q6[16]}}, q6[16:6]};
             q7 <= q6 - {{6{i6[16]}}, i6[16:6]};
          end
        else
          begin
             a7 <= a6[12:0] - 13'd2607;
             i7 <= i6 - {{6{q6[16]}}, q6[16:6]};
             q7 <= q6 + {{6{i6[16]}}, i6[16:6]};
          end // else: !if(a6[14])
        /* 0.448 degrees */
        if(a7[12])
          begin
             a8 <= a7[11:0] + 12'd1304;
             i8 <= i7 + {{7{q7[16]}}, q7[16:7]};
             q8 <= q7 - {{7{i7[16]}}, i7[16:7]};
          end
        else
          begin
             a8 <= a7[11:0] - 12'd1304;
             i8<= i7 - {{7{q7[16]}}, q7[16:7]};
             q8 <= q7 + {{7{i7[16]}}, i7[16:7]};
          end // else: !if(a7[14])
        /* 0.224 degrees */
        if(a8[11])
          begin
             a9 <= a8[10:0] + 11'd652;
             i9 <= i8 + {{8{q8[16]}}, q8[16:8]};
             q9 <= q8 - {{8{i8[16]}}, i8[16:8]};
          end
        else
          begin
             a9 <= a8[10:0] - 11'd652;
             i9 <= i8 - {{8{q8[16]}}, q8[16:8]};
             q9 <= q8 + {{8{i8[16]}}, i8[16:8]};
          end // else: !if(a8[11])
        /* 0.1119 degrees */
        if(a9[10])
          begin
             a10 <= a9[9:0] + 10'd326;
             i10 <= i9 + {{9{q9[16]}}, q9[16:9]};
             q10 <= q9 - {{9{i9[16]}}, i9[16:9]};
          end
        else
          begin
             a10 <= a9[9:0] - 10'd326;
             i10 <= i9 - {{9{q9[16]}}, q9[16:9]};
             q10 <= q9 + {{9{i9[16]}}, i9[16:9]};
          end // else: !if(a9[10])
        /* 0.05595 degrees */
        if(a10[9])
          begin
             a11 <= a10[8:0] + 9'd163;
             i11 <= i10 + {{10{q10[16]}}, q10[16:10]};
             q11 <= q10 - {{10{i10[16]}}, i10[16:10]};
          end
        else
          begin
             a11 <= a10[8:0] - 9'd163;
             i11 <= i10 - {{10{q10[16]}}, q10[16:10]};
             q11 <= q10 + {{10{i10[16]}}, i10[16:10]};
          end // else: !if(a10[9])
        /* 0.02798 degrees */
        if(a11[8])
          begin
             a12 <= a11[7:0] + 8'd81;
             i12 <= i11 + {{11{q11[16]}}, q11[16:11]};
             q12 <= q11 - {{11{i11[16]}}, i11[16:11]};
          end
        else
          begin
             a12 <= a11[7:0] - 8'd81;
             i12 <= i11 - {{11{q11[16]}}, q11[16:11]};
             q12 <= q11 + {{11{i11[16]}}, i11[16:11]};
          end // else: !if(a11[8])
        /* 0.01399 degrees */
        if(a12[7])
          begin
             a13 <= a12[6:0] + 7'd41;
             i13 <= i12 + {{12{q12[16]}}, q12[16:12]};
             q13 <= q12 - {{12{i12[16]}}, i12[16:12]};
          end
        else
          begin
             a13 <= a12[6:0] - 7'd41;
             i13 <= i12 - {{12{q12[16]}}, q12[16:12]};
             q13 <= q12 + {{12{i12[16]}}, i12[16:12]};
          end // else: !if(a12[7])
        /* 0.00699 degrees */
        if(a13[6])
          begin 
             a14 <= a13[5:0] + 6'd20;
             i14 <= i13 + {{13{q13[16]}}, q13[16:13]};
             q14 <= q13 - {{13{i13[16]}}, i13[16:13]};
          end
        else
          begin
             a14 <= a13[5:0] - 6'd20;
             i14 <= i13 - {{13{q13[16]}}, q13[16:13]};
             q14 <= q13 + {{13{i13[16]}}, i13[16:13]};
          end // else: !if(a13[6])
        /* 0.00350 degrees */
        if(a14[5])
          begin
             a15 <= a14[4:0] + 5'd10;
             i15 <= i14 + {{14{q14[16]}}, q14[16:14]};
             q15 <= q14 - {{14{i14[16]}}, i14[16:14]};
          end
        else
          begin
             a15 <= a14[4:0] - 5'd10;
             i15 <= i14 - {{14{q14[16]}}, q14[16:14]};
             q15 <= q14 + {{14{i14[16]}}, i14[16:14]};
          end // else: !if(a14[5])
        /* 0.00175 degrees */
        if(a15[4])
          begin
             i16 <= i15 + {{15{q15[16]}}, q15[16:15]};
             q16 <= q15 - {{15{i15[16]}}, i15[16:15]};
          end
        else
          begin
             i16 <= i15 - {{15{q15[16]}}, q15[16:15]};
             q16 <= q15 + {{15{i15[16]}}, i15[16:15]};
          end // else: !if(a15[4])      
     end // always @ (posedge clk)
   assign iout = i16;
   assign qout = q16;
endmodule //cordic
