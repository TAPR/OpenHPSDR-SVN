// Copyright (c) 2007 Christopher T. Day (AE6VK@Yahoo.com)
//
// HPSDR - High Performance Software Defined Radio
//
// Interface between Janus OnBoard discrete hardware and the
// JanusCPLD system.
// 
// The software supports the Alpha1 version of the Janus board.
//
//
// This program is free software; you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation; either version 2 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA 
// 02111-1307  USA
//
//
module OnBoard_interface (
	// Pins
	input	OnBoard_XO_out,
	output	OnBoard_PWMFilter_I,
	output	OnBoard_PWMFilter_Q,
	input	OnBoard_PTT,
	inout	OnBoard_J7Header1,
	inout	OnBoard_J7Header2,
	inout	OnBoard_J7Header3,
	inout	OnBoard_J7Header4,
	// Wires
	output	Clk,
	input	PWMI,
	input	PWMQ,
	output	PTT,
	inout	[3:0] TestHeader
	);
	
	// Assemble the full interface from its components.	
	XO_interface XO (OnBoard_XO_out, Clk);
	
	PWMFilter_interface PWMFilter (OnBoard_PWMFilter_I, 
								   OnBoard_PWMFilter_Q,
								   PWMI, PWMQ);
		
	PTT_interface PTTHrdw (OnBoard_PTT, PTT);
	
	TestHeader_interface TestHeaderJ7 (OnBoard_J7Header1,
									   OnBoard_J7Header2,
									   OnBoard_J7Header3,
									   OnBoard_J7Header4,
									   TestHeader);

endmodule
