module cROM(clk, addr, data, reset);

	input clk;
	input [7:0] addr;
	input reset;
	output signed [23:0] data;

	reg [23:0] data;

	always @(posedge clk) begin
		if (reset)
			data <= 0;
		else begin
			case(addr)
				8'd0: data <= 24'sh0;
				8'd1: data <= 24'sha;
				8'd2: data <= 24'sh14;
				8'd3: data <= 24'sh1e;
				8'd4: data <= 24'sh28;
				8'd5: data <= 24'sh32;
				8'd6: data <= 24'sh3c;
				8'd7: data <= 24'sh46;
				8'd8: data <= 24'sh50;
				8'd9: data <= 24'sh5a;
				8'd10: data <= 24'sh64;
				8'd11: data <= 24'sh6e;
				8'd12: data <= 24'sh78;
				8'd13: data <= 24'sh82;
				8'd14: data <= 24'sh8c;
				8'd15: data <= 24'sh96;
				8'd16: data <= 24'sha0;
				8'd17: data <= 24'shaa;
				8'd18: data <= 24'shb4;
				8'd19: data <= 24'shbe;
				8'd20: data <= 24'shc8;
				8'd21: data <= 24'shd2;
				8'd22: data <= 24'shdc;
				8'd23: data <= 24'she6;
				8'd24: data <= 24'shf0;
				8'd25: data <= 24'shfa;
				8'd26: data <= 24'sh104;
				8'd27: data <= 24'sh10e;
				8'd28: data <= 24'sh118;
				8'd29: data <= 24'sh122;
				8'd30: data <= 24'sh12c;
				8'd31: data <= 24'sh136;
				8'd32: data <= 24'sh140;
				8'd33: data <= 24'sh14a;
				8'd34: data <= 24'sh154;
				8'd35: data <= 24'sh15e;
				8'd36: data <= 24'sh168;
				8'd37: data <= 24'sh172;
				8'd38: data <= 24'sh17c;
				8'd39: data <= 24'sh186;
				8'd40: data <= 24'sh190;
				8'd41: data <= 24'sh19a;
				8'd42: data <= 24'sh1a4;
				8'd43: data <= 24'sh1ae;
				8'd44: data <= 24'sh1b8;
				8'd45: data <= 24'sh1c2;
				8'd46: data <= 24'sh1cc;
				8'd47: data <= 24'sh1d6;
				8'd48: data <= 24'sh1e0;
				8'd49: data <= 24'sh1ea;
				8'd50: data <= 24'sh1f4;
				8'd51: data <= 24'sh1fe;
				8'd52: data <= 24'sh208;
				8'd53: data <= 24'sh212;
				8'd54: data <= 24'sh21c;
				8'd55: data <= 24'sh226;
				8'd56: data <= 24'sh230;
				8'd57: data <= 24'sh23a;
				8'd58: data <= 24'sh244;
				8'd59: data <= 24'sh24e;
				8'd60: data <= 24'sh258;
				8'd61: data <= 24'sh262;
				8'd62: data <= 24'sh26c;
				8'd63: data <= 24'sh276;
				8'd64: data <= 24'sh280;
				8'd65: data <= 24'sh28a;
				8'd66: data <= 24'sh294;
				8'd67: data <= 24'sh29e;
				8'd68: data <= 24'sh2a8;
				8'd69: data <= 24'sh2b2;
				8'd70: data <= 24'sh2bc;
				8'd71: data <= 24'sh2c6;
				8'd72: data <= 24'sh2d0;
				8'd73: data <= 24'sh2da;
				8'd74: data <= 24'sh2e4;
				8'd75: data <= 24'sh2ee;
				8'd76: data <= 24'sh2f8;
				8'd77: data <= 24'sh302;
				8'd78: data <= 24'sh30c;
				8'd79: data <= 24'sh316;
				8'd80: data <= 24'sh320;
				8'd81: data <= 24'sh32a;
				8'd82: data <= 24'sh334;
				8'd83: data <= 24'sh33e;
				8'd84: data <= 24'sh348;
				8'd85: data <= 24'sh352;
				8'd86: data <= 24'sh35c;
				8'd87: data <= 24'sh366;
				8'd88: data <= 24'sh370;
				8'd89: data <= 24'sh37a;
				8'd90: data <= 24'sh384;
				8'd91: data <= 24'sh38e;
				8'd92: data <= 24'sh398;
				8'd93: data <= 24'sh3a2;
				8'd94: data <= 24'sh3ac;
				8'd95: data <= 24'sh3b6;
				8'd96: data <= 24'sh3c0;
				8'd97: data <= 24'sh3ca;
				8'd98: data <= 24'sh3d4;
				8'd99: data <= 24'sh3de;
				8'd100: data <= 24'sh3e8;
				8'd101: data <= 24'sh3f2;
				8'd102: data <= 24'sh3fc;
				8'd103: data <= 24'sh406;
				8'd104: data <= 24'sh410;
				8'd105: data <= 24'sh41a;
				8'd106: data <= 24'sh424;
				8'd107: data <= 24'sh42e;
				8'd108: data <= 24'sh438;
				8'd109: data <= 24'sh442;
				8'd110: data <= 24'sh44c;
				8'd111: data <= 24'sh456;
				8'd112: data <= 24'sh460;
				8'd113: data <= 24'sh46a;
				8'd114: data <= 24'sh474;
				8'd115: data <= 24'sh47e;
				8'd116: data <= 24'sh488;
				8'd117: data <= 24'sh492;
				8'd118: data <= 24'sh49c;
				8'd119: data <= 24'sh4a6;
				8'd120: data <= 24'sh4b0;
				8'd121: data <= 24'sh4ba;
				8'd122: data <= 24'sh4c4;
				8'd123: data <= 24'sh4ce;
				8'd124: data <= 24'sh4d8;
				8'd125: data <= 24'sh4e2;
				8'd126: data <= 24'sh4ec;
				8'd127: data <= 24'sh4f6;
				8'd128: data <= 24'sh500;
				8'd129: data <= 24'sh50a;
				8'd130: data <= 24'sh514;
				8'd131: data <= 24'sh51e;
				8'd132: data <= 24'sh528;
				8'd133: data <= 24'sh532;
				8'd134: data <= 24'sh53c;
				8'd135: data <= 24'sh546;
				8'd136: data <= 24'sh550;
				8'd137: data <= 24'sh55a;
				8'd138: data <= 24'sh564;
				8'd139: data <= 24'sh56e;
				8'd140: data <= 24'sh578;
				8'd141: data <= 24'sh582;
				8'd142: data <= 24'sh58c;
				8'd143: data <= 24'sh596;
				8'd144: data <= 24'sh5a0;
				8'd145: data <= 24'sh5aa;
				8'd146: data <= 24'sh5b4;
				8'd147: data <= 24'sh5be;
				8'd148: data <= 24'sh5c8;
				8'd149: data <= 24'sh5d2;
				8'd150: data <= 24'sh5dc;
				8'd151: data <= 24'sh5e6;
				8'd152: data <= 24'sh5f0;
				8'd153: data <= 24'sh5fa;
				8'd154: data <= 24'sh604;
				8'd155: data <= 24'sh60e;
				8'd156: data <= 24'sh618;
				8'd157: data <= 24'sh622;
				8'd158: data <= 24'sh62c;
				8'd159: data <= 24'sh636;
				8'd160: data <= 24'sh640;
				8'd161: data <= 24'sh64a;
				8'd162: data <= 24'sh654;
				8'd163: data <= 24'sh65e;
				8'd164: data <= 24'sh668;
				8'd165: data <= 24'sh672;
				8'd166: data <= 24'sh67c;
				8'd167: data <= 24'sh686;
				8'd168: data <= 24'sh690;
				8'd169: data <= 24'sh69a;
				8'd170: data <= 24'sh6a4;
				8'd171: data <= 24'sh6ae;
				8'd172: data <= 24'sh6b8;
				8'd173: data <= 24'sh6c2;
				8'd174: data <= 24'sh6cc;
				8'd175: data <= 24'sh6d6;
				8'd176: data <= 24'sh6e0;
				8'd177: data <= 24'sh6ea;
				8'd178: data <= 24'sh6f4;
				8'd179: data <= 24'sh6fe;
				8'd180: data <= 24'sh708;
				8'd181: data <= 24'sh712;
				8'd182: data <= 24'sh71c;
				8'd183: data <= 24'sh726;
				8'd184: data <= 24'sh730;
				8'd185: data <= 24'sh73a;
				8'd186: data <= 24'sh744;
				8'd187: data <= 24'sh74e;
				8'd188: data <= 24'sh758;
				8'd189: data <= 24'sh762;
				8'd190: data <= 24'sh76c;
				8'd191: data <= 24'sh776;
				8'd192: data <= 24'sh780;
				8'd193: data <= 24'sh78a;
				8'd194: data <= 24'sh794;
				8'd195: data <= 24'sh79e;
				8'd196: data <= 24'sh7a8;
				8'd197: data <= 24'sh7b2;
				8'd198: data <= 24'sh7bc;
				8'd199: data <= 24'sh7c6;
				8'd200: data <= 24'sh7d0;
				8'd201: data <= 24'sh7da;
				8'd202: data <= 24'sh7e4;
				8'd203: data <= 24'sh7ee;
				8'd204: data <= 24'sh7f8;
				8'd205: data <= 24'sh802;
				8'd206: data <= 24'sh80c;
				8'd207: data <= 24'sh816;
				8'd208: data <= 24'sh820;
				8'd209: data <= 24'sh82a;
				8'd210: data <= 24'sh834;
				8'd211: data <= 24'sh83e;
				8'd212: data <= 24'sh848;
				8'd213: data <= 24'sh852;
				8'd214: data <= 24'sh85c;
				8'd215: data <= 24'sh866;
				8'd216: data <= 24'sh870;
				8'd217: data <= 24'sh87a;
				8'd218: data <= 24'sh884;
				8'd219: data <= 24'sh88e;
				8'd220: data <= 24'sh898;
				8'd221: data <= 24'sh8a2;
				8'd222: data <= 24'sh8ac;
				8'd223: data <= 24'sh8b6;
				8'd224: data <= 24'sh8c0;
				8'd225: data <= 24'sh8ca;
				8'd226: data <= 24'sh8d4;
				8'd227: data <= 24'sh8de;
				8'd228: data <= 24'sh8e8;
				8'd229: data <= 24'sh8f2;
				8'd230: data <= 24'sh8fc;
				8'd231: data <= 24'sh906;
				8'd232: data <= 24'sh910;
				8'd233: data <= 24'sh91a;
				8'd234: data <= 24'sh924;
				8'd235: data <= 24'sh92e;
				8'd236: data <= 24'sh938;
				8'd237: data <= 24'sh942;
				8'd238: data <= 24'sh94c;
				8'd239: data <= 24'sh956;
				8'd240: data <= 24'sh960;
				8'd241: data <= 24'sh96a;
				8'd242: data <= 24'sh974;
				8'd243: data <= 24'sh97e;
				8'd244: data <= 24'sh988;
				8'd245: data <= 24'sh992;
				8'd246: data <= 24'sh99c;
				8'd247: data <= 24'sh9a6;
				8'd248: data <= 24'sh9b0;
				8'd249: data <= 24'sh9ba;
				8'd250: data <= 24'sh9c4;
				8'd251: data <= 24'sh9ce;
				8'd252: data <= 24'sh9d8;
				8'd253: data <= 24'sh9e2;
				8'd254: data <= 24'sh9ec;
				8'd255: data <= 24'sh9f6;
				default: data <= 24'sh0;
			endcase
		end
	end

endmodule
